module dataMem(
	input logic [7:0] addr,
	input logic [7:0] write_data,
	input logic mem_write,
	input logic mem_read,
	output logic [7:0] data_out
);

//fill in guts
	logic[7:0] Core[256];
	
	always_comb begin 
	//do this later
	end

endmodule